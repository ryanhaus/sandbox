module top(
    input clk,
    input rst,

    output hsync,
    output vsync,
    output [7:0] red,
    output [7:0] green,
    output [7:0] blue
);

endmodule
