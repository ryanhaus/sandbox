module tca9539();

endmodule
